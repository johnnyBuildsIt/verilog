module uart_rx
#(parameter CLKS_PER_BIT = 217)(
  input        i_Clock,
  input        i_RX_Serial,
  output       o_RX_DV,
  output [7:0] o_RX_Byte
);



endmodule