module seven_seg_test (
  output o_Segment1_A,
  output o_Segment1_B,
  output o_Segment1_C,
  output o_Segment1_D,
  output o_Segment1_E,
  output o_Segment1_F,
  output o_Segment1_G);

assign o_Segment1_A = 1'b0;
assign o_Segment1_B = 1'b1;
assign o_Segment1_C = 1'b0;
assign o_Segment1_D = 1'b0;
assign o_Segment1_E = 1'b1;
assign o_Segment1_F = 1'b0;
assign o_Segment1_G = 1'b0;
    
endmodule